library IEEE;
use IEEE.std_logic_1164.all;

entity Lab_3_1_1131417 is
    port(
        CLK : in std_logic;
        DIN : in std_logic;
        Q   : out std_logic_vector(7 downto 0)
    );
end Lab_3_1_1131417;

architecture RDL of Lab_3_1_1131417 is
    signal reg : std_logic_vector(7 downto 0);
begin
    process(CLK)
    begin
        if rising_edge(CLK) then
            reg <= reg(6 downto 0) & DIN; -- �����ADIN �i S0
        end if;
    end process;
    Q <= reg;
end RDL;

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_Lab_3_1_1131417 is
end tb_Lab_3_1_1131417;

architecture sim of tb_Lab_3_1_1131417 is
    signal CLK : std_logic := '0';
    signal DIN : std_logic := '0';
    signal Q   : std_logic_vector(7 downto 0);
begin
    -- DUT
    uut: entity work.Lab_3_1_1131417
        port map(CLK => CLK, DIN => DIN, Q => Q);

    -- Clock 10ns
    CLK <= not CLK after 5 ns;

    -- DIN 20ns
    process
    begin
        DIN <= '1'; wait for 20 ns;
        DIN <= '0'; wait for 20 ns;
        DIN <= '1'; wait for 20 ns;
        DIN <= '1'; wait for 20 ns;
        DIN <= '0'; wait for 20 ns;
        DIN <= '1'; wait for 20 ns;
        wait;
    end process;
end sim;