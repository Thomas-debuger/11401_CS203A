library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity minsec_timer is
    generic(
        CLK_FREQ : integer := 50000000
    );
    port (
        clk   : in  std_logic;
        hex0  : out std_logic_vector(7 downto 0); -- ��Ӧ�
        hex1  : out std_logic_vector(7 downto 0); -- ��Q�� + �p���I
        hex2  : out std_logic_vector(7 downto 0); -- ���Ӧ�
        hex3  : out std_logic_vector(7 downto 0)  -- ���Q��
    );
end minsec_timer;

architecture rtl of minsec_timer is

    -- BCD �p�ɭ�
    signal m_tens  : integer range 0 to 5 := 5;
    signal m_units : integer range 0 to 9 := 9;
    signal s_tens  : integer range 0 to 5 := 5;
    signal s_units : integer range 0 to 9 := 7;

    -- 1Hz tick
    constant COUNT_1HZ : integer := CLK_FREQ - 1;
    signal cnt_1hz  : integer := 0;
    signal tick_1hz : std_logic := '0';

    -- BCD �� 7�q�]active-low�Adp = �̥��� bit�^
    function bcd7seg(x : integer; dp : std_logic) return std_logic_vector is
        variable seg : std_logic_vector(7 downto 0);
    begin
        case x is
            when 0 => seg := dp & "1000000";
            when 1 => seg := dp & "1111001";
            when 2 => seg := dp & "0100100";
            when 3 => seg := dp & "0110000";
            when 4 => seg := dp & "0011001";
            when 5 => seg := dp & "0010010";
            when 6 => seg := dp & "0000010";
            when 7 => seg := dp & "1111000";
            when 8 => seg := dp & "0000000";
            when 9 => seg := dp & "0010000";
            when others => seg := dp & "1111111";
        end case;
        return seg;
    end function;

begin

    -------------------------------------------------------------
    -- 1Hz tick
    -------------------------------------------------------------
    process(clk)
    begin
        if rising_edge(clk) then
            if cnt_1hz = COUNT_1HZ then
                cnt_1hz  <= 0;
                tick_1hz <= '1';
            else
                cnt_1hz  <= cnt_1hz + 1;
                tick_1hz <= '0';
            end if;
        end if;
    end process;

    -------------------------------------------------------------
    -- ����p�ɾ�
    -------------------------------------------------------------
    process(clk)
    begin
        if rising_edge(clk) then
            if tick_1hz = '1' then

                if s_units < 9 then
                    s_units <= s_units + 1;
                else
                    s_units <= 0;

                    if s_tens < 5 then
                        s_tens <= s_tens + 1;
                    else
                        s_tens <= 0;

                        if m_units < 9 then
                            m_units <= m_units + 1;
                        else
                            m_units <= 0;

                            if m_tens < 5 then
                                m_tens <= m_tens + 1;
                            else
                                m_tens <= 0;
                            end if;
                        end if;

                    end if;

                end if;

            end if;
        end if;
    end process;

    -------------------------------------------------------------
    -- ��X�C�q�]�p���I�b HEX1�^
    -- dp = 0 �G, 1 �� (active-low)
    -------------------------------------------------------------
    hex0 <= bcd7seg(s_units, '1'); -- no dp
    hex1 <= bcd7seg(s_tens, '1'); -- dp ON (�b��Ʀr����)
    hex2 <= bcd7seg(m_units, '0');
    hex3 <= bcd7seg(m_tens, '1');

end rtl;